module testbench;
    test_ifu IFU();
endmodule
